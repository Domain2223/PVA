magic
tech scmos
timestamp 1714630292
<< metal1 >>
rect 579 820 1181 824
rect 571 812 1173 816
rect 563 804 1165 808
rect 555 796 1157 800
rect 547 788 1149 792
rect 539 780 1141 784
rect 531 772 1133 776
rect 523 764 1125 768
rect 1123 697 1181 701
rect 757 680 764 684
rect 445 656 765 660
rect 1123 589 1173 593
rect 511 567 644 571
rect 749 567 753 571
rect 763 563 767 576
rect 579 559 646 563
rect 753 559 767 563
rect 383 533 408 537
rect 423 533 451 537
rect 417 502 459 506
rect 463 502 467 506
rect 471 502 475 506
rect 479 502 483 506
rect 487 502 491 506
rect 495 502 499 506
rect 503 502 507 506
rect 383 481 408 485
rect 753 479 757 559
rect 1123 481 1165 485
rect 503 475 636 479
rect 749 475 757 479
rect 571 467 638 471
rect 753 464 764 468
rect 394 395 409 399
rect 753 387 757 464
rect 495 383 628 387
rect 749 383 757 387
rect 563 375 630 379
rect 1123 373 1157 377
rect 753 356 765 360
rect -4 301 0 305
rect -12 293 -8 297
rect 753 295 757 356
rect 487 291 620 295
rect 749 291 757 295
rect -20 285 -16 289
rect 555 283 622 287
rect -28 277 -24 281
rect 1123 265 1149 269
rect 384 261 407 265
rect 447 263 584 265
rect 447 261 588 263
rect 580 259 588 261
rect 753 248 764 252
rect 441 234 445 235
rect -46 229 -42 233
rect 384 209 407 213
rect 447 211 584 213
rect 447 209 588 211
rect 580 207 588 209
rect 753 203 757 248
rect 479 199 612 203
rect 749 199 757 203
rect 547 191 614 195
rect 1123 156 1141 160
rect 753 139 763 143
rect 753 111 757 139
rect 471 107 604 111
rect 749 107 757 111
rect 539 99 606 103
rect 753 55 764 59
rect 753 27 757 55
rect 1123 48 1133 52
rect 398 22 425 26
rect 749 23 757 27
rect 763 19 767 35
rect 463 15 596 19
rect 749 15 767 19
rect 531 7 598 11
rect 756 -1 764 3
rect 756 -13 760 -1
rect 610 -17 614 -13
rect 749 -17 760 -13
rect -77 -56 -72 -52
rect 1123 -60 1125 -56
rect -77 -64 -72 -60
rect 455 -77 588 -73
rect 749 -77 763 -73
rect 523 -85 590 -81
rect 186 -109 921 -105
rect 222 -117 957 -113
<< m2contact >>
rect 575 820 579 824
rect 1181 820 1185 824
rect 567 812 571 816
rect 1173 812 1177 816
rect 559 804 563 808
rect 1165 804 1169 808
rect 551 796 555 800
rect 1157 796 1161 800
rect 543 788 547 792
rect 1149 788 1153 792
rect 535 780 539 784
rect 1141 780 1145 784
rect 527 772 531 776
rect 1133 772 1137 776
rect 519 764 523 768
rect 1125 764 1129 768
rect 1181 697 1185 701
rect 753 680 757 684
rect 441 656 445 660
rect 765 656 769 660
rect -81 598 -77 602
rect 1173 589 1177 593
rect 507 567 511 571
rect 753 567 757 571
rect 575 559 579 563
rect 451 533 455 537
rect 409 501 413 505
rect 459 502 463 506
rect 467 502 471 506
rect 475 502 479 506
rect 483 502 487 506
rect 491 502 495 506
rect 499 502 503 506
rect 507 502 511 506
rect 1165 481 1169 485
rect 499 475 503 479
rect 567 467 571 471
rect 409 395 413 399
rect 491 383 495 387
rect 559 375 563 379
rect 1157 373 1161 377
rect 483 291 487 295
rect 551 283 555 287
rect 1149 265 1153 269
rect -71 229 -67 233
rect 409 229 413 233
rect 425 229 429 233
rect 441 230 445 234
rect 475 199 479 203
rect 543 191 547 195
rect 1141 156 1145 160
rect -48 128 -44 132
rect 467 107 471 111
rect -81 100 -77 104
rect 535 99 539 103
rect 1133 48 1137 52
rect 425 22 429 26
rect 459 15 463 19
rect 527 7 531 11
rect 1125 -60 1129 -56
rect 610 -69 614 -65
rect 451 -77 455 -73
rect 519 -85 523 -81
rect 182 -109 186 -105
rect 921 -109 925 -105
rect 218 -117 222 -113
rect 957 -117 961 -113
<< metal2 >>
rect -81 104 -77 598
rect -71 233 -67 477
rect 106 208 110 376
rect 114 261 118 429
rect 182 277 186 421
rect 218 269 222 413
rect 409 399 413 501
rect 409 233 413 395
rect 441 234 445 656
rect 394 192 398 199
rect 386 127 390 134
rect 378 29 382 36
rect 425 26 429 229
rect 182 -105 186 -52
rect 218 -113 222 -64
rect 342 -67 346 -60
rect 451 -73 455 533
rect 507 506 511 567
rect 459 19 463 502
rect 467 111 471 502
rect 475 203 479 502
rect 483 295 487 502
rect 491 387 495 502
rect 499 479 503 502
rect 519 -81 523 764
rect 527 11 531 772
rect 535 103 539 780
rect 543 195 547 788
rect 551 287 555 796
rect 559 379 563 804
rect 567 471 571 812
rect 575 563 579 820
rect 753 571 757 680
rect 610 -41 614 -37
rect 1125 -56 1129 764
rect 921 -105 925 -97
rect 957 -113 961 -98
rect 1125 -101 1129 -60
rect 1133 52 1137 772
rect 1133 -101 1137 48
rect 1141 160 1145 780
rect 1141 -101 1145 156
rect 1149 269 1153 788
rect 1149 -101 1153 265
rect 1157 377 1161 796
rect 1157 -101 1161 373
rect 1165 485 1169 804
rect 1165 -101 1169 481
rect 1173 593 1177 812
rect 1173 -101 1177 589
rect 1181 701 1185 820
rect 1181 -101 1185 697
use 8BitAdder  8BitAdder_0
timestamp 1714603105
transform 1 0 588 0 1 -69
box -6 -32 165 706
use INV  INV_0
timestamp 1711561836
transform 1 0 407 0 1 481
box -4 0 20 59
use OR2  OR2_0
timestamp 1712274593
transform 1 0 407 0 1 209
box -6 0 44 62
use RegEn8  RegEn8_0
timestamp 1714615249
transform 1 0 763 0 1 -53
box -4 -48 366 825
use RotationDetector  RotationDetector_0
timestamp 1714588023
transform 1 0 0 0 1 0
box -77 -96 398 277
use RotationDetector  RotationDetector_1
timestamp 1714588023
transform 1 0 0 0 1 373
box -77 -96 398 277
<< labels >>
rlabel metal2 1127 -99 1127 -99 1 Q0
rlabel metal2 1135 -99 1135 -99 1 Q1
rlabel metal2 1143 -99 1143 -99 1 Q2
rlabel metal2 1151 -99 1151 -99 1 Q3
rlabel metal2 1159 -99 1159 -99 1 Q4
rlabel metal2 1167 -99 1167 -99 1 Q5
rlabel metal2 1175 -99 1175 -99 1 Q6
rlabel metal1 -76 -54 -76 -54 3 RST
rlabel metal1 -76 -62 -76 -62 3 CLK
rlabel metal2 108 347 108 347 1 VSS
rlabel metal2 117 345 117 345 1 VDD
rlabel metal2 411 459 411 459 1 rot1
rlabel metal1 439 504 439 504 1 rot1`
rlabel metal2 427 167 427 167 1 rot2
rlabel metal2 443 288 443 288 1 en
rlabel metal2 396 196 396 196 1 q2
rlabel metal2 388 131 388 131 1 q2b
rlabel metal2 379 34 379 34 1 q1
rlabel metal2 344 -64 344 -64 1 q1b
rlabel metal1 -44 231 -44 231 1 r2r`
rlabel m2contact -46 130 -46 130 1 r2in`
rlabel metal1 -26 279 -26 279 1 s1
rlabel metal1 -18 287 -18 287 1 s1`
rlabel metal1 -11 295 -11 295 1 s2
rlabel metal1 -2 303 -2 303 1 s2`
rlabel metal1 757 -75 757 -74 1 a0
rlabel metal1 756 17 756 17 1 a1
rlabel metal1 753 109 753 109 1 a2
rlabel metal1 755 201 755 201 1 a3
rlabel metal1 754 293 754 293 1 a4
rlabel metal1 755 407 755 407 1 a5
rlabel metal1 755 494 755 494 1 a6
rlabel metal2 755 614 755 614 1 a7
rlabel metal2 1183 -99 1183 -99 7 Q7
rlabel metal2 -69 341 -69 341 1 fwd
rlabel metal2 -79 340 -79 340 3 bwd
<< end >>
