magic
tech scmos
timestamp 1711596499
use INV  INV_0 ~/cmpe480-s24/PVA
timestamp 1711561836
transform 1 0 4 0 1 -1
box -4 0 20 59
use NAND2  NAND2_0
timestamp 1711563584
transform 1 0 20 0 1 -1
box -6 0 34 62
<< labels >>
rlabel polycontact 8 17 8 17 1 A
rlabel polycontact 35 27 35 27 1 B
rlabel metal1 44 27 44 27 1 Y
rlabel metal1 8 53 8 53 1 VDD
rlabel metal1 8 1 8 1 1 VSS
<< end >>
