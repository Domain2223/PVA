magic
tech scmos
timestamp 1711488442
<< metal1 >>
rect 0 52 150 56
rect 138 32 142 36
rect 34 24 38 28
rect 70 24 74 28
rect 106 24 110 28
rect 174 24 182 28
rect 210 24 214 28
rect 0 0 6 4
rect 26 -8 110 -4
rect 114 -8 138 -4
rect 182 -8 210 -4
rect 38 -16 66 -12
rect 70 -16 166 -12
rect 62 -24 130 -20
rect 134 -24 202 -20
rect 78 -32 94 -28
rect 106 -32 218 -28
<< m2contact >>
rect 2 48 6 52
rect 146 48 150 52
rect 22 32 26 36
rect 34 32 38 36
rect 58 32 62 36
rect 70 32 74 36
rect 94 32 98 36
rect 106 32 110 36
rect 130 32 134 36
rect 166 32 170 36
rect 178 32 182 36
rect 202 32 206 36
rect 214 32 218 36
rect 2 28 6 32
rect 146 28 150 32
rect 138 24 142 28
rect 66 20 70 24
rect 102 20 106 24
rect 210 20 214 24
rect 22 -8 26 -4
rect 110 -8 114 -4
rect 138 -8 142 -4
rect 178 -8 182 -4
rect 210 -8 214 -4
rect 34 -16 38 -12
rect 66 -16 70 -12
rect 166 -16 170 -12
rect 58 -24 62 -20
rect 130 -24 134 -20
rect 202 -24 206 -20
rect 74 -32 78 -28
rect 94 -32 98 -28
rect 102 -32 106 -28
rect 218 -32 222 -28
<< metal2 >>
rect 2 32 6 48
rect 22 -4 26 32
rect 34 -12 38 32
rect 58 -20 62 32
rect 66 -12 70 20
rect 74 -28 78 36
rect 94 -28 98 32
rect 102 -28 106 20
rect 110 -4 114 36
rect 130 -20 134 32
rect 146 32 150 48
rect 138 -4 142 24
rect 166 -12 170 32
rect 178 -4 182 32
rect 202 -20 206 32
rect 210 -4 214 20
rect 218 -28 222 36
use NAND3  NAND3_0
timestamp 1709762292
transform 1 0 0 0 1 0
box -6 0 42 62
use NAND3  NAND3_1
timestamp 1709762292
transform 1 0 36 0 1 0
box -6 0 42 62
use NAND3  NAND3_2
timestamp 1709762292
transform 1 0 72 0 1 0
box -6 0 42 62
use NAND3  NAND3_3
timestamp 1709762292
transform 1 0 108 0 1 0
box -6 0 42 62
use NAND3  NAND3_4
timestamp 1709762292
transform 1 0 144 0 1 0
box -6 0 42 62
use NAND3  NAND3_5
timestamp 1709762292
transform 1 0 180 0 1 0
box -6 0 42 62
<< labels >>
rlabel metal1 140 34 140 34 1 D
rlabel metal1 4 54 4 54 1 VDD
rlabel metal1 4 2 4 2 1 VSS
rlabel m2contact 76 -30 76 -30 1 CLK
rlabel metal1 176 26 176 26 1 Q
rlabel metal1 212 26 212 26 1 Qb
rlabel m2contact 60 -22 60 -22 1 RS
<< end >>
