magic
tech scmos
timestamp 1711561843
<< nwell >>
rect -6 42 34 66
<< ntransistor >>
rect 8 8 10 12
rect 18 8 20 12
<< ptransistor >>
rect 8 48 10 52
rect 18 48 20 52
<< ndiffusion >>
rect 7 8 8 12
rect 10 8 18 12
rect 20 8 22 12
<< pdiffusion >>
rect 6 48 8 52
rect 10 48 12 52
rect 16 48 18 52
rect 20 48 22 52
<< ndcontact >>
rect 3 8 7 12
rect 22 8 26 12
<< pdcontact >>
rect 2 48 6 52
rect 12 48 16 52
rect 22 48 26 52
<< psubstratepcontact >>
rect 3 0 7 4
<< nsubstratencontact >>
rect 2 56 6 60
<< polysilicon >>
rect 8 52 10 54
rect 18 52 20 54
rect 8 30 10 48
rect 18 30 20 48
rect 7 26 10 30
rect 17 26 20 30
rect 8 12 10 26
rect 18 12 20 26
rect 8 6 10 8
rect 18 6 20 8
<< polycontact >>
rect 3 26 7 30
rect 13 26 17 30
<< metal1 >>
rect 0 56 2 60
rect 6 56 28 60
rect 2 52 6 56
rect 22 52 26 56
rect 12 44 16 48
rect 12 40 26 44
rect 22 12 26 40
rect 3 4 7 8
rect 0 0 3 4
rect 7 0 26 4
<< labels >>
rlabel psubstratepcontact 5 2 5 2 1 VSS
rlabel nsubstratencontact 4 58 4 58 1 VDD
rlabel polycontact 5 28 5 28 1 A
rlabel polycontact 15 28 15 28 1 B
rlabel metal1 24 28 24 28 1 Y
<< end >>
