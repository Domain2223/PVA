magic
tech scmos
timestamp 1711563584
<< nwell >>
rect -6 38 34 62
<< ntransistor >>
rect 8 8 10 12
rect 18 8 20 12
<< ptransistor >>
rect 8 44 10 48
rect 18 44 20 48
<< ndiffusion >>
rect 7 8 8 12
rect 10 8 18 12
rect 20 8 22 12
<< pdiffusion >>
rect 6 44 8 48
rect 10 44 12 48
rect 16 44 18 48
rect 20 44 22 48
<< ndcontact >>
rect 3 8 7 12
rect 22 8 26 12
<< pdcontact >>
rect 2 44 6 48
rect 12 44 16 48
rect 22 44 26 48
<< psubstratepcontact >>
rect 3 0 7 4
<< nsubstratencontact >>
rect 2 52 6 56
<< polysilicon >>
rect 8 48 10 50
rect 18 48 20 50
rect 8 30 10 44
rect 18 30 20 44
rect 7 26 10 30
rect 17 26 20 30
rect 8 12 10 26
rect 18 12 20 26
rect 8 6 10 8
rect 18 6 20 8
<< polycontact >>
rect 3 26 7 30
rect 13 26 17 30
<< metal1 >>
rect 0 52 2 56
rect 6 52 28 56
rect 2 48 6 52
rect 22 48 26 52
rect 12 40 16 44
rect 12 36 26 40
rect 22 12 26 36
rect 3 4 7 8
rect 0 0 3 4
rect 7 0 28 4
<< labels >>
rlabel psubstratepcontact 5 2 5 2 1 VSS
rlabel polycontact 5 28 5 28 1 A
rlabel polycontact 15 28 15 28 1 B
rlabel metal1 24 28 24 28 1 Y
rlabel nsubstratencontact 4 54 4 54 1 VDD
<< end >>
