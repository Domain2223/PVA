magic
tech scmos
timestamp 1710799370
<< nwell >>
rect -4 38 20 63
<< ntransistor >>
rect 7 8 9 12
<< ptransistor >>
rect 7 44 9 52
<< ndiffusion >>
rect 6 8 7 12
rect 9 8 10 12
<< pdiffusion >>
rect 6 44 7 52
rect 9 44 10 52
<< ndcontact >>
rect 2 8 6 12
rect 10 8 14 12
<< pdcontact >>
rect 2 44 6 52
rect 10 44 14 52
<< psubstratepcontact >>
rect 6 0 10 4
<< nsubstratencontact >>
rect 6 56 10 60
<< polysilicon >>
rect 7 52 9 54
rect 7 20 9 44
rect 6 16 9 20
rect 7 12 9 16
rect 7 6 9 8
<< polycontact >>
rect 2 16 6 20
<< metal1 >>
rect 0 56 6 60
rect 10 56 16 60
rect 2 52 6 56
rect 10 12 14 44
rect 2 4 6 8
rect 0 0 6 4
rect 10 0 16 4
<< labels >>
rlabel metal1 4 2 4 2 1 VSS
rlabel polycontact 4 18 4 18 1 A
rlabel metal1 12 18 12 18 1 Y
rlabel metal1 4 58 4 58 1 VDD
<< end >>
