magic
tech scmos
timestamp 1711591893
<< nwell >>
rect -4 38 54 62
<< ntransistor >>
rect 8 8 10 12
rect 18 8 20 12
rect 28 8 30 12
rect 38 8 40 12
<< ptransistor >>
rect 8 44 10 48
rect 18 44 20 48
rect 28 44 30 48
rect 38 44 40 48
<< ndiffusion >>
rect 6 8 8 12
rect 10 8 18 12
rect 20 8 28 12
rect 30 8 38 12
rect 40 8 42 12
<< pdiffusion >>
rect 6 44 8 48
rect 10 44 12 48
rect 16 44 18 48
rect 20 44 22 48
rect 26 44 28 48
rect 30 44 32 48
rect 36 44 38 48
rect 40 44 42 48
<< ndcontact >>
rect 2 8 6 12
rect 42 8 46 12
<< pdcontact >>
rect 2 44 6 48
rect 12 44 16 48
rect 22 44 26 48
rect 32 44 36 48
rect 42 44 46 48
<< psubstratepcontact >>
rect 2 0 6 4
<< nsubstratencontact >>
rect 2 52 6 56
<< polysilicon >>
rect 8 48 10 50
rect 18 48 20 50
rect 28 48 30 50
rect 38 48 40 50
rect 8 32 10 44
rect 7 28 10 32
rect 8 12 10 28
rect 18 24 20 44
rect 28 32 30 44
rect 27 28 30 32
rect 17 20 20 24
rect 18 12 20 20
rect 28 12 30 28
rect 38 24 40 44
rect 37 20 40 24
rect 38 12 40 20
rect 8 6 10 8
rect 18 6 20 8
rect 28 6 30 8
rect 38 6 40 8
<< polycontact >>
rect 3 28 7 32
rect 23 28 27 32
rect 13 20 17 24
rect 33 20 37 24
<< metal1 >>
rect 0 52 2 56
rect 6 52 48 56
rect 12 48 16 52
rect 32 48 36 52
rect 2 40 6 44
rect 22 40 26 44
rect 42 40 46 44
rect 2 36 46 40
rect 42 12 46 36
rect 2 4 6 8
rect 0 0 2 4
rect 6 0 48 4
<< labels >>
rlabel polycontact 5 30 5 30 1 A
rlabel polycontact 15 22 15 22 1 B
rlabel polycontact 25 30 25 30 1 C
rlabel polycontact 35 22 35 22 1 D
rlabel metal1 8 2 8 2 1 VSS
rlabel metal1 8 54 8 54 1 VDD
rlabel metal1 44 24 44 24 1 Y
<< end >>
