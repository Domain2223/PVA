magic
tech scmos
timestamp 1714632880
<< metal1 >>
rect 1213 731 1374 735
rect 1221 679 1374 683
rect 1124 663 1209 667
rect 1124 611 1217 615
rect 1221 611 1223 615
rect 503 479 587 483
rect 901 479 963 483
rect 591 443 663 447
rect 871 443 897 447
rect 503 427 595 431
rect 909 427 963 431
rect 599 391 663 395
rect 879 391 905 395
rect 1134 120 1270 124
rect 1130 112 1138 116
rect 1142 112 1250 116
rect 1254 112 1268 116
rect 1130 104 1146 108
rect 1150 104 1242 108
rect 1246 104 1268 108
rect 1130 96 1154 100
rect 1158 96 1234 100
rect 1238 96 1268 100
rect 1130 88 1162 92
rect 1166 88 1226 92
rect 1230 88 1268 92
rect 1130 80 1170 84
rect 1174 80 1218 84
rect 1222 80 1268 84
rect 1130 72 1178 76
rect 1182 72 1210 76
rect 1214 72 1268 76
rect 1130 64 1186 68
rect 1190 64 1202 68
rect 1206 64 1268 68
rect 609 36 662 40
rect 1258 28 1270 32
rect 609 24 621 28
rect 617 12 621 24
rect 666 23 713 27
rect 1266 16 1396 20
rect -5 -20 56 -16
rect 60 -20 677 -16
rect 681 -20 1388 -16
rect 1392 -20 1606 -16
rect 268 -44 617 -40
rect 276 -52 597 -48
rect 284 -60 589 -56
rect 292 -68 581 -64
rect -20 -130 1290 -126
rect 1294 -130 1350 -126
rect -20 -138 1298 -134
rect 1302 -138 1350 -134
rect -20 -146 1306 -142
rect 1310 -146 1350 -142
rect -20 -154 1314 -150
rect 1318 -154 1350 -150
rect -20 -162 1322 -158
rect 1326 -162 1350 -158
rect -20 -170 1330 -166
rect 1334 -170 1350 -166
rect -20 -178 1338 -174
rect 1342 -178 1350 -174
rect -20 -186 1346 -182
<< m2contact >>
rect 1209 731 1213 735
rect 1217 679 1221 683
rect 1209 663 1213 667
rect 1217 611 1221 615
rect 587 479 591 483
rect 897 479 901 483
rect 587 443 591 447
rect 897 443 901 447
rect 595 427 599 431
rect 905 427 909 431
rect 595 391 599 395
rect 905 391 909 395
rect 1130 120 1134 124
rect 1270 120 1274 124
rect 1138 112 1142 116
rect 1250 112 1254 116
rect 1146 104 1150 108
rect 1242 104 1246 108
rect 1154 96 1158 100
rect 1234 96 1238 100
rect 1162 88 1166 92
rect 1226 88 1230 92
rect 1170 80 1174 84
rect 1218 80 1222 84
rect 1396 79 1400 83
rect 1178 72 1182 76
rect 1210 72 1214 76
rect 1186 64 1190 68
rect 1202 64 1206 68
rect 662 36 666 40
rect 581 28 585 32
rect 589 28 593 32
rect 597 28 601 32
rect 1202 28 1206 32
rect 1210 28 1214 32
rect 1218 28 1222 32
rect 1226 28 1230 32
rect 1234 28 1238 32
rect 1242 28 1246 32
rect 1250 28 1254 32
rect 1270 28 1274 32
rect 662 23 666 27
rect 713 23 717 27
rect 1396 16 1400 20
rect 617 8 621 12
rect 56 -20 60 -16
rect 677 -20 681 -16
rect 1388 -20 1392 -16
rect 264 -44 268 -40
rect 617 -44 621 -40
rect 272 -52 276 -48
rect 597 -52 601 -48
rect 280 -60 284 -56
rect 589 -60 593 -56
rect 288 -68 292 -64
rect 581 -68 585 -64
rect 1290 -130 1294 -126
rect 1298 -138 1302 -134
rect 1306 -146 1310 -142
rect 1314 -154 1318 -150
rect 1322 -162 1326 -158
rect 1330 -170 1334 -166
rect 1338 -178 1342 -174
rect 1346 -186 1350 -182
<< metal2 >>
rect 1209 667 1213 731
rect 1209 487 1213 663
rect 1217 615 1221 679
rect 1217 487 1221 611
rect 587 447 591 479
rect 897 447 901 479
rect 595 395 599 427
rect 905 395 909 427
rect 1202 68 1206 124
rect 56 -16 60 27
rect 92 23 96 27
rect 264 -40 268 0
rect 272 -48 276 0
rect 280 -56 284 0
rect 288 -64 292 0
rect 581 -64 585 28
rect 589 -56 593 28
rect 597 -48 601 28
rect 662 27 666 36
rect 1202 32 1206 64
rect 1210 76 1214 124
rect 1210 32 1214 72
rect 1218 84 1222 124
rect 1218 32 1222 80
rect 1226 92 1230 124
rect 1226 32 1230 88
rect 1234 100 1238 124
rect 1234 32 1238 96
rect 1242 108 1246 124
rect 1242 32 1246 104
rect 1250 116 1254 124
rect 1250 32 1254 112
rect 1270 32 1274 120
rect 662 21 666 23
rect 617 -40 621 8
rect 677 -16 681 27
rect 1290 -126 1294 53
rect 1290 -186 1294 -130
rect 1298 -134 1302 53
rect 1298 -186 1302 -138
rect 1306 -142 1310 53
rect 1306 -186 1310 -146
rect 1314 -150 1318 53
rect 1314 -186 1318 -154
rect 1322 -158 1326 53
rect 1322 -186 1326 -162
rect 1330 -166 1334 53
rect 1330 -186 1334 -170
rect 1338 -174 1342 53
rect 1338 -186 1342 -178
rect 1346 -182 1350 53
rect 1388 -16 1392 71
rect 1396 20 1400 79
rect 2596 9 2600 825
rect 2604 9 2608 61
rect 2612 9 2616 61
rect 2620 9 2624 61
rect 2628 9 2632 61
rect 2636 9 2640 61
rect 2644 9 2648 61
rect 2652 9 2656 61
use COUNTER4  COUNTER4_1
timestamp 1714614791
transform 1 0 36 0 1 27
box -36 -27 533 777
use COUNTER4  COUNTER4_2
timestamp 1714614791
transform 1 0 657 0 1 27
box -36 -27 533 777
use DELTAX  DELTAX_0
timestamp 1714632880
transform 1 0 1368 0 1 99
box -78 -99 1288 992
use NOR4  NOR4_0
timestamp 1711564571
transform 1 0 575 0 1 0
box -6 0 46 62
use NOR8  NOR8_0
timestamp 1711565688
transform 1 0 1196 0 1 0
box -6 0 78 62
<< labels >>
rlabel metal2 94 25 94 25 1 CLK
rlabel metal1 -3 -18 -3 -18 1 RST
rlabel metal1 -18 -184 -18 -184 2 A0
rlabel metal1 -18 -176 -18 -176 3 A1
rlabel metal1 -18 -168 -18 -168 3 A2
rlabel metal1 -18 -160 -18 -160 3 A3
rlabel metal1 -18 -152 -18 -152 3 A4
rlabel metal1 -18 -144 -18 -144 3 A5
rlabel metal1 -18 -136 -18 -136 3 A6
rlabel metal1 -17 -128 -17 -128 3 A7
rlabel metal2 2654 11 2654 11 7 Y0
rlabel metal2 2646 11 2646 11 1 Y1
rlabel metal2 2638 11 2638 11 1 Y2
rlabel metal2 2630 11 2630 11 1 Y3
rlabel metal2 2622 11 2622 11 1 Y4
rlabel metal2 2614 11 2614 11 1 Y5
rlabel metal2 2606 11 2606 11 1 Y6
rlabel metal2 2598 11 2598 11 1 Y7
rlabel m2contact 589 481 589 481 1 VDD
<< end >>
