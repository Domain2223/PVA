magic
tech scmos
timestamp 1711561836
<< nwell >>
rect -4 34 20 59
<< ntransistor >>
rect 7 8 9 12
<< ptransistor >>
rect 7 40 9 48
<< ndiffusion >>
rect 6 8 7 12
rect 9 8 10 12
<< pdiffusion >>
rect 6 40 7 48
rect 9 40 10 48
<< ndcontact >>
rect 2 8 6 12
rect 10 8 14 12
<< pdcontact >>
rect 2 40 6 48
rect 10 40 14 48
<< psubstratepcontact >>
rect 6 0 10 4
<< nsubstratencontact >>
rect 6 52 10 56
<< polysilicon >>
rect 7 48 9 50
rect 7 20 9 40
rect 6 16 9 20
rect 7 12 9 16
rect 7 6 9 8
<< polycontact >>
rect 2 16 6 20
<< metal1 >>
rect 0 52 6 56
rect 10 52 16 56
rect 2 48 6 52
rect 10 12 14 40
rect 2 4 6 8
rect 0 0 6 4
rect 10 0 16 4
<< labels >>
rlabel metal1 4 2 4 2 1 VSS
rlabel polycontact 4 18 4 18 1 A
rlabel metal1 12 18 12 18 1 Y
rlabel metal1 4 54 4 54 1 VDD
<< end >>
