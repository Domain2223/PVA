magic
tech scmos
timestamp 1714589065
<< nwell >>
rect 158 52 161 56
<< metal1 >>
rect -35 696 0 700
rect -37 656 -33 660
rect -35 644 0 648
rect -29 636 0 640
rect 3 636 6 640
rect 161 636 163 640
rect 11 628 14 632
rect 161 628 163 632
rect 123 620 127 624
rect -35 604 0 608
rect -37 564 -33 568
rect -35 552 0 556
rect -29 544 1 548
rect 4 544 6 548
rect 161 544 164 548
rect 11 536 14 540
rect 131 536 161 540
rect 123 528 127 532
rect -35 512 0 516
rect -37 472 -33 476
rect -35 460 0 464
rect -29 452 0 456
rect 3 452 6 456
rect 161 452 163 456
rect 11 444 14 448
rect 131 444 161 448
rect 123 436 127 440
rect -35 420 0 424
rect -37 380 -33 384
rect -36 368 1 372
rect -29 360 0 364
rect 3 360 6 364
rect 161 360 163 364
rect 11 352 14 356
rect 131 352 161 356
rect 123 344 127 348
rect -35 328 0 332
rect -37 288 -33 292
rect -35 276 0 280
rect -29 268 0 272
rect 4 268 6 272
rect 161 268 163 272
rect 12 260 14 264
rect 131 260 161 264
rect 123 252 127 256
rect -36 236 0 240
rect -38 196 -34 200
rect -36 184 0 188
rect -30 176 0 180
rect 3 176 6 180
rect 161 176 163 180
rect 12 168 14 172
rect 131 168 161 172
rect 123 160 127 164
rect -36 144 0 148
rect -38 104 -34 108
rect -36 92 0 96
rect -30 84 0 88
rect 4 84 6 88
rect 161 84 163 88
rect 12 76 14 80
rect 131 76 161 80
rect 123 68 127 72
rect -36 52 0 56
rect 158 52 161 56
rect -38 12 -34 16
rect -36 0 0 4
rect 161 0 163 4
rect -30 -8 0 -4
rect 161 -8 163 -4
rect 131 -16 155 -12
rect 161 -16 163 -12
<< m2contact >>
rect 54 696 58 700
rect -33 656 -29 660
rect 94 644 98 648
rect -33 636 -29 640
rect 127 620 131 624
rect 54 604 58 608
rect -33 564 -29 568
rect 94 552 98 556
rect -33 544 -29 548
rect 127 536 131 540
rect 127 528 131 532
rect 54 512 58 516
rect -33 472 -29 476
rect 94 460 98 464
rect -33 452 -29 456
rect 127 444 131 448
rect 127 436 131 440
rect 54 420 58 424
rect -33 380 -29 384
rect 94 368 98 372
rect -33 360 -29 364
rect 127 352 131 356
rect 127 344 131 348
rect 54 328 58 332
rect -33 288 -29 292
rect 94 276 98 280
rect -33 268 -29 272
rect 127 260 131 264
rect 127 252 131 256
rect 54 236 58 240
rect -34 196 -30 200
rect 94 184 98 188
rect -34 176 -30 180
rect 127 168 131 172
rect 127 160 131 164
rect 54 144 58 148
rect -34 104 -30 108
rect 94 92 98 96
rect -34 84 -30 88
rect 127 76 131 80
rect 127 68 131 72
rect 54 52 58 56
rect -34 12 -30 16
rect 94 0 98 4
rect -34 -8 -30 -4
rect 127 -16 131 -12
<< metal2 >>
rect -33 640 -29 656
rect 54 608 58 696
rect -33 548 -29 564
rect 54 516 58 604
rect -33 456 -29 472
rect 54 424 58 512
rect -33 364 -29 380
rect 54 332 58 420
rect -33 272 -29 288
rect 54 240 58 328
rect -34 180 -30 196
rect 54 148 58 236
rect -34 88 -30 104
rect 54 56 58 144
rect 94 556 98 644
rect 94 464 98 552
rect 127 540 131 620
rect 94 372 98 460
rect 127 448 131 528
rect 94 280 98 368
rect 127 356 131 436
rect 94 188 98 276
rect 127 264 131 344
rect 94 96 98 184
rect 127 172 131 252
rect -34 -4 -30 12
rect 94 4 98 92
rect 127 80 131 160
rect 127 -12 131 68
use FullAdder  FullAdder_0
timestamp 1713982514
transform 1 0 0 0 1 0
box -6 -32 165 62
use FullAdder  FullAdder_1
timestamp 1713982514
transform 1 0 0 0 1 92
box -6 -32 165 62
use FullAdder  FullAdder_2
timestamp 1713982514
transform 1 0 0 0 1 184
box -6 -32 165 62
use FullAdder  FullAdder_3
timestamp 1713982514
transform 1 0 0 0 1 276
box -6 -32 165 62
use FullAdder  FullAdder_4
timestamp 1713982514
transform 1 0 0 0 1 368
box -6 -32 165 62
use FullAdder  FullAdder_5
timestamp 1713982514
transform 1 0 0 0 1 460
box -6 -32 165 62
use FullAdder  FullAdder_6
timestamp 1713982514
transform 1 0 0 0 1 552
box -6 -32 165 62
use FullAdder  FullAdder_7
timestamp 1713982514
transform 1 0 0 0 1 644
box -6 -32 165 62
use XOR2  XOR2_0
timestamp 1711599452
transform 1 0 -156 0 1 0
box 0 -24 126 62
use XOR2  XOR2_1
timestamp 1711599452
transform 1 0 -152 0 1 -97
box 0 -24 126 62
use XOR2  XOR2_2
timestamp 1711599452
transform 1 0 -156 0 1 184
box 0 -24 126 62
use XOR2  XOR2_3
timestamp 1711599452
transform 1 0 -156 0 1 92
box 0 -24 126 62
use XOR2  XOR2_4
timestamp 1711599452
transform 1 0 -155 0 1 276
box 0 -24 126 62
use XOR2  XOR2_5
timestamp 1711599452
transform 1 0 -155 0 1 368
box 0 -24 126 62
use XOR2  XOR2_6
timestamp 1711599452
transform 1 0 -155 0 1 460
box 0 -24 126 62
use XOR2  XOR2_7
timestamp 1711599452
transform 1 0 -155 0 1 552
box 0 -24 126 62
use XOR2  XOR2_8
timestamp 1711599452
transform 1 0 -155 0 1 644
box 0 -24 126 62
<< labels >>
rlabel metal1 162 -6 162 -6 1 S0
rlabel metal1 5 86 5 86 1 A1
rlabel metal1 13 78 13 78 1 B1
rlabel metal1 162 86 162 86 1 S1
rlabel metal1 5 178 5 178 1 A2
rlabel metal1 13 170 13 170 1 B2
rlabel metal1 162 178 162 178 1 S2
rlabel metal1 5 270 5 270 1 A3
rlabel metal1 13 262 13 262 1 B3
rlabel metal1 162 270 162 270 1 S3
rlabel metal1 5 362 5 362 1 A4
rlabel metal1 12 354 12 354 1 B4
rlabel metal1 162 362 162 362 1 S4
rlabel metal1 5 454 5 454 1 A5
rlabel metal1 12 446 12 446 1 B5
rlabel metal1 162 454 162 454 1 S5
rlabel metal1 5 546 5 546 1 A6
rlabel metal1 13 538 13 538 1 B6
rlabel metal1 162 546 162 546 1 S6
rlabel metal1 5 638 5 638 1 A7
rlabel metal1 12 630 12 630 1 B7
rlabel metal1 162 638 162 638 1 S7
rlabel metal1 162 630 162 630 1 Cout
rlabel metal1 162 2 162 2 1 VSS
rlabel metal1 159 54 159 54 1 VDD
<< end >>
