magic
tech scmos
timestamp 1711593671
<< metal1 >>
rect 0 52 6 56
rect 30 24 46 28
rect 102 24 118 28
rect 178 24 190 28
rect 0 0 6 4
rect 26 -8 66 -4
rect 70 -8 150 -4
rect 170 -7 210 -3
rect 6 -16 14 -12
rect 18 -16 86 -12
rect 90 -16 158 -12
rect 178 -16 214 -12
rect 6 -24 50 -20
rect 54 -24 78 -20
rect 98 -24 138 -20
rect 34 -32 122 -28
rect 62 -40 102 -36
rect 106 -40 194 -36
<< m2contact >>
rect 130 52 134 56
rect 202 52 206 56
rect 174 24 178 28
rect 6 20 10 24
rect 14 20 18 24
rect 22 20 26 24
rect 30 20 34 24
rect 50 20 54 24
rect 58 20 62 24
rect 66 20 70 24
rect 78 20 82 24
rect 86 20 90 24
rect 94 20 98 24
rect 102 20 106 24
rect 122 20 126 24
rect 130 20 134 24
rect 138 20 142 24
rect 150 20 154 24
rect 158 20 162 24
rect 166 20 170 24
rect 194 20 198 24
rect 202 20 206 24
rect 210 20 214 24
rect 6 -8 10 -4
rect 22 -8 26 -4
rect 66 -8 70 -4
rect 150 -8 154 -4
rect 166 -7 170 -3
rect 210 -7 214 -3
rect 14 -16 18 -12
rect 86 -16 90 -12
rect 158 -16 162 -12
rect 174 -16 178 -12
rect 50 -24 54 -20
rect 78 -24 82 -20
rect 94 -24 98 -20
rect 138 -24 142 -20
rect 30 -32 34 -28
rect 122 -32 126 -28
rect 58 -40 62 -36
rect 102 -40 106 -36
rect 194 -40 198 -36
<< metal2 >>
rect 130 24 134 52
rect 202 24 206 52
rect 6 -4 10 20
rect 14 -12 18 20
rect 22 -4 26 20
rect 30 -28 34 20
rect 50 -20 54 20
rect 58 -36 62 20
rect 66 -4 70 20
rect 78 -20 82 20
rect 86 -12 90 20
rect 94 -20 98 20
rect 102 -36 106 20
rect 122 -28 126 20
rect 138 -20 142 20
rect 150 -4 154 20
rect 158 -12 162 20
rect 166 -3 170 20
rect 174 -12 178 24
rect 194 -36 198 20
rect 210 -3 214 20
use NAND3  NAND3_0
timestamp 1711593430
transform 1 0 0 0 1 0
box -6 0 42 62
use NAND3  NAND3_1
timestamp 1711593430
transform 1 0 36 0 1 0
box -6 0 42 62
use NAND3  NAND3_2
timestamp 1711593430
transform 1 0 72 0 1 0
box -6 0 42 62
use NAND3  NAND3_3
timestamp 1711593430
transform 1 0 108 0 1 0
box -6 0 42 62
use NAND3  NAND3_4
timestamp 1711593430
transform 1 0 144 0 1 0
box -6 0 42 62
use NAND3  NAND3_5
timestamp 1711593430
transform 1 0 180 0 1 0
box -6 0 42 62
<< labels >>
rlabel m2contact 8 -6 8 -6 1 D
rlabel m2contact 16 -14 16 -14 1 RST
rlabel m2contact 52 -22 52 -22 1 CLK
rlabel metal1 4 2 4 2 1 VSS
rlabel metal1 4 54 4 54 1 VDD
rlabel m2contact 212 -5 212 -5 1 Q
rlabel metal1 213 -14 213 -14 1 Qb
<< end >>
